library verilog;
use verilog.vl_types.all;
entity Simple_vlg_vec_tst is
end Simple_vlg_vec_tst;
