library verilog;
use verilog.vl_types.all;
entity lab15_part2_vlg_vec_tst is
end lab15_part2_vlg_vec_tst;
